module first(a,b,c);
input a,b;
output c;
assign c=a&b;
endmodule


// module first(a, b);

// input a;
// output b;
// assign b =~a;

// endmodule